entity test is port( a, b, c : in bit;
                     z : out bit); end test;

architecture data_flow of test is
begin
end data_flow;
